`define VX_ADDRESS 1
