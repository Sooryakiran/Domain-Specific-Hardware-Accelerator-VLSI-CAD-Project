// Defines the address of the memory mapped Vector Accelerator
`define VX_ADDRESS 1
