`define VX_NEG 1
`define VX_REDUCE_MIN 11
