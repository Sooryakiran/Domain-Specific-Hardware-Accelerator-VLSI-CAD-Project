`define WORD_LENGTH 32
`define DATA_LENGTH 32
`define PC_SIZE 32

`define SMALL_WIDTH True